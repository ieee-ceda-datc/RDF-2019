MACRO AND2x11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x11_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.412 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.412 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.496 2.952 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.664 0.444 2.736 0.636 ; 
    END 
  END A
END AND2x11_ASAP7_75t_SL

MACRO AND2x13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x13_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.844 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.844 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.496 3.384 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.096 0.444 3.168 0.636 ; 
    END 
  END A
END AND2x13_ASAP7_75t_SL

MACRO AND2x14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x14_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 3.060 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 3.060 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.528 0.496 3.600 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.444 3.384 0.636 ; 
    END 
  END A
END AND2x14_ASAP7_75t_SL

MACRO AND2x3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x3_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.684 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.496 1.224 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.444 1.008 0.636 ; 
    END 
  END A
END AND2x3_ASAP7_75t_SL

MACRO AND2x4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x4_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.008 0.180 ; 
        RECT 0.936 0.180 1.008 0.900 ; 
        RECT 0.396 0.900 1.008 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.496 1.440 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.444 1.224 0.636 ; 
    END 
  END A
END AND2x4_ASAP7_75t_SL

MACRO AND2x6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x6_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.440 0.180 ; 
        RECT 1.368 0.180 1.440 0.900 ; 
        RECT 0.396 0.900 1.440 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.496 1.872 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.444 1.656 0.636 ; 
    END 
  END A
END AND2x6_ASAP7_75t_SL

MACRO AND2x7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x7_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.548 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.548 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.496 2.088 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.444 1.872 0.636 ; 
    END 
  END A
END AND2x7_ASAP7_75t_SL

MACRO AND2x9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x9_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.980 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.980 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.496 2.520 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.444 2.304 0.636 ; 
    END 
  END A
END AND2x9_ASAP7_75t_SL

MACRO AO221x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO221x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END C
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END A2
END AO221x1_ASAP7_75t_SL

MACRO AO222x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO222x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.468 0.180 ; 
        RECT 0.288 0.180 0.360 0.756 ; 
        RECT 0.360 0.684 0.468 0.756 ; 
    END 
  END Y
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END C2
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B2
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END B1
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END C1
END AO222x2_ASAP7_75t_SL

MACRO AO332x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO332x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.444 0.792 0.636 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.444 0.576 0.636 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.444 1.008 0.636 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.444 1.224 0.636 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.444 1.440 0.636 ; 
    END 
  END B2
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.444 1.656 0.636 ; 
    END 
  END B3
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.444 1.872 0.636 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.444 2.088 0.636 ; 
    END 
  END C1
END AO332x1_ASAP7_75t_SL

MACRO AOI21x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.324 1.440 0.396 ; 
        RECT 0.720 0.396 0.792 0.576 ; 
        RECT 1.368 0.396 1.440 0.576 ; 
    END 
  END A2
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END B
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A1
END AOI21x1_ASAP7_75t_SL

MACRO AOI22x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.180 1.548 0.252 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
        RECT 0.144 0.684 0.900 0.756 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 1.008 0.396 ; 
        RECT 0.288 0.396 0.360 0.576 ; 
        RECT 0.936 0.396 1.008 0.576 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.324 1.872 0.396 ; 
        RECT 1.152 0.396 1.224 0.576 ; 
        RECT 1.800 0.396 1.872 0.576 ; 
    END 
  END B1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END A2
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.348 0.504 1.460 0.576 ; 
    END 
  END B2
END AOI22x1_ASAP7_75t_SL

MACRO AOI322xp5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI322xp5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END B1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END C1
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END C2
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.252 1.872 0.324 ; 
        RECT 1.800 0.324 1.872 0.756 ; 
        RECT 1.476 0.756 1.872 0.828 ; 
    END 
  END Y
END AOI322xp5_ASAP7_75t_SL

MACRO AOI332xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI332xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 1.332 0.324 ; 
        RECT 0.072 0.324 0.144 0.828 ; 
        RECT 0.144 0.756 0.468 0.828 ; 
    END 
  END Y
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A1
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B3
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END A3
END AOI332xp33_ASAP7_75t_SL

MACRO AOI333xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI333xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 1.548 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN C3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END C3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A1
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END C1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A3
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B3
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B1
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C2
END AOI333xp33_ASAP7_75t_SL

MACRO BUFx11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx11_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.412 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.412 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.664 0.424 2.736 0.656 ; 
    END 
  END A
END BUFx11_ASAP7_75t_SL

MACRO BUFx12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx12_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 2.628 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 2.628 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.424 2.952 0.656 ; 
    END 
  END A
END BUFx12_ASAP7_75t_SL

MACRO BUFx14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx14_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 3.060 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 3.060 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.424 3.384 0.656 ; 
    END 
  END A
END BUFx14_ASAP7_75t_SL

MACRO BUFx15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx15_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 3.276 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 3.276 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.528 0.424 3.600 0.656 ; 
    END 
  END A
END BUFx15_ASAP7_75t_SL

MACRO BUFx4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx4_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.900 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 0.900 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A
END BUFx4_ASAP7_75t_SL

MACRO BUFx5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.116 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.116 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A
END BUFx5_ASAP7_75t_SL

MACRO BUFx8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx8_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.872 0.180 ; 
        RECT 1.800 0.180 1.872 0.900 ; 
        RECT 0.396 0.900 1.872 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.996 0.504 2.108 0.576 ; 
    END 
  END A
END BUFx8_ASAP7_75t_SL

MACRO DFFHQNx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx1_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.484 0.360 0.596 ; 
    END 
  END CLK
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.484 1.224 0.596 ; 
    END 
  END D
  PIN QN
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.852 0.324 4.248 0.396 ; 
        RECT 4.176 0.396 4.248 0.684 ; 
        RECT 3.852 0.684 4.248 0.756 ; 
    END 
  END QN
END DFFHQNx1_ASAP7_75t_SL

MACRO DHLx2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx2_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.324 3.168 0.396 ; 
        RECT 3.096 0.396 3.168 0.684 ; 
        RECT 2.988 0.684 3.168 0.756 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx2_ASAP7_75t_SL

MACRO DHLx3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx3_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.108 3.492 0.180 ; 
        RECT 2.880 0.180 2.952 0.972 ; 
        RECT 2.952 0.900 3.492 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx3_ASAP7_75t_SL

MACRO DHLx5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx5_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.108 4.032 0.180 ; 
        RECT 3.960 0.180 4.032 0.900 ; 
        RECT 2.988 0.900 4.032 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx5_ASAP7_75t_SL

MACRO DHLx6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx6_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.108 4.032 0.180 ; 
        RECT 3.960 0.180 4.032 0.900 ; 
        RECT 2.988 0.900 4.032 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx6_ASAP7_75t_SL

MACRO FAx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FAx1_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN CON
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.160 0.756 0.704 0.828 ; 
    END 
  END CON
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.348 0.252 2.324 0.324 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.376 0.612 2.756 0.684 ; 
    END 
  END A
  PIN CI
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.396 2.540 0.468 ; 
    END 
  END CI
  PIN SN
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.888 0.108 2.864 0.180 ; 
    END 
  END SN
END FAx1_ASAP7_75t_SL

MACRO INVx11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx11_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.736 0.180 ; 
        RECT 2.664 0.180 2.736 0.900 ; 
        RECT 0.396 0.900 2.736 0.972 ; 
    END 
  END Y
END INVx11_ASAP7_75t_SL

MACRO INVx12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx12_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.736 0.180 ; 
        RECT 2.664 0.180 2.736 0.900 ; 
        RECT 0.396 0.900 2.736 0.972 ; 
    END 
  END Y
END INVx12_ASAP7_75t_SL

MACRO INVx14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx14_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.168 0.180 ; 
        RECT 3.096 0.180 3.168 0.900 ; 
        RECT 0.396 0.900 3.168 0.972 ; 
    END 
  END Y
END INVx14_ASAP7_75t_SL

MACRO INVx16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx16_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.600 0.180 ; 
        RECT 3.528 0.180 3.600 0.900 ; 
        RECT 0.396 0.900 3.600 0.972 ; 
    END 
  END Y
END INVx16_ASAP7_75t_SL

MACRO INVx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx1_ASAP7_75t_SL 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.252 0.576 0.324 ; 
        RECT 0.504 0.324 0.576 0.756 ; 
        RECT 0.396 0.756 0.576 0.828 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
END INVx1_ASAP7_75t_SL

MACRO INVx2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx2_ASAP7_75t_SL 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.324 0.576 0.396 ; 
        RECT 0.504 0.396 0.576 0.684 ; 
        RECT 0.396 0.684 0.576 0.756 ; 
    END 
  END Y
END INVx2_ASAP7_75t_SL

MACRO INVx3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx3_ASAP7_75t_SL 0 0 ; 
  SIZE 1.080 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.684 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
END INVx3_ASAP7_75t_SL

MACRO INVx5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.116 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.116 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.504 1.008 0.576 ; 
    END 
  END A
END INVx5_ASAP7_75t_SL

MACRO INVx6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx6_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.504 1.008 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 1.332 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 1.332 0.972 ; 
    END 
  END Y
END INVx6_ASAP7_75t_SL

MACRO 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN  0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.108 3.492 0.180 ; 
        RECT 2.880 0.180 2.952 0.972 ; 
        RECT 2.952 0.900 3.492 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END 

MACRO INVx9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx9_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.304 0.180 ; 
        RECT 2.232 0.180 2.304 0.900 ; 
        RECT 0.396 0.900 2.304 0.972 ; 
    END 
  END Y
END INVx9_ASAP7_75t_SL

MACRO NAND2x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.468 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.900 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END B
END NAND2x1_ASAP7_75t_SL

MACRO NOR4xp25_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR4xp25_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.900 0.180 ; 
        RECT 0.072 0.180 0.144 0.828 ; 
        RECT 0.144 0.756 0.252 0.828 ; 
    END 
  END Y
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
END NOR4xp25_ASAP7_75t_SL

MACRO NOR5xp2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR5xp2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.116 0.180 ; 
        RECT 0.072 0.180 0.144 0.828 ; 
        RECT 0.144 0.756 0.252 0.828 ; 
    END 
  END Y
  PIN E
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END E
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
END NOR5xp2_ASAP7_75t_SL

MACRO OA33x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA33x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A2
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B3
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END B1
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.288 0.396 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
END OA33x2_ASAP7_75t_SL

MACRO OAI21xp5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.080 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.684 0.324 ; 
        RECT 0.072 0.324 0.144 0.828 ; 
        RECT 0.144 0.756 0.468 0.828 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END B
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
END OAI21xp5_ASAP7_75t_SL

MACRO OAI22xp5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI22xp5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.828 0.252 1.224 0.324 ; 
        RECT 1.152 0.324 1.224 0.756 ; 
        RECT 0.612 0.756 1.224 0.828 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B2
END OAI22xp5_ASAP7_75t_SL

MACRO OAI321xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI321xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.260 0.252 1.656 0.324 ; 
        RECT 1.584 0.324 1.656 0.900 ; 
        RECT 0.828 0.900 1.656 0.972 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B2
END OAI321xp33_ASAP7_75t_SL

MACRO OAI322xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI322xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.468 0.324 ; 
        RECT 0.072 0.324 0.144 0.828 ; 
        RECT 0.144 0.756 1.332 0.828 ; 
    END 
  END Y
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B2
END OAI322xp33_ASAP7_75t_SL

MACRO OAI32xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI32xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.044 0.252 1.440 0.324 ; 
        RECT 1.368 0.324 1.440 0.756 ; 
        RECT 0.828 0.756 1.440 0.828 ; 
    END 
  END Y
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
END OAI32xp33_ASAP7_75t_SL

MACRO OAI331xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI331xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.072 0.324 0.144 0.828 ; 
        RECT 0.144 0.756 1.116 0.828 ; 
    END 
  END Y
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B3
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A3
END OAI331xp33_ASAP7_75t_SL

MACRO OAI333xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI333xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.684 0.180 ; 
        RECT 0.072 0.180 0.144 0.828 ; 
        RECT 0.144 0.756 1.548 0.828 ; 
    END 
  END Y
  PIN C3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END C3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A1
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END C1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A3
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B3
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B1
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C2
END OAI333xp33_ASAP7_75t_SL

MACRO OR2x10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x10_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.304 0.180 ; 
        RECT 2.232 0.180 2.304 0.900 ; 
        RECT 0.396 0.900 2.304 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.664 0.424 2.736 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END A
END OR2x10_ASAP7_75t_SL

MACRO OR2x11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x11_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.412 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.412 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.424 2.952 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.664 0.424 2.736 0.656 ; 
    END 
  END A
END OR2x11_ASAP7_75t_SL

MACRO OR2x12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x12_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.736 0.180 ; 
        RECT 2.664 0.180 2.736 0.900 ; 
        RECT 0.396 0.900 2.736 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.096 0.424 3.168 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.424 2.952 0.656 ; 
    END 
  END A
END OR2x12_ASAP7_75t_SL

MACRO OR2x13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x13_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.844 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.844 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.424 3.384 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.096 0.424 3.168 0.656 ; 
    END 
  END A
END OR2x13_ASAP7_75t_SL

MACRO OR2x15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x15_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 3.276 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 3.276 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.744 0.424 3.816 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.528 0.424 3.600 0.656 ; 
    END 
  END A
END OR2x15_ASAP7_75t_SL

MACRO OR2x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.468 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A
END OR2x2_ASAP7_75t_SL

MACRO OR2x3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x3_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.684 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A
END OR2x3_ASAP7_75t_SL

MACRO OR4x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR4x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
END OR4x1_ASAP7_75t_SL

MACRO XNOR2x10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x10_ASAP7_75t_SL 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 2.412 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 3.060 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.724 0.504 3.836 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.644 0.504 2.756 0.576 ; 
    END 
  END B
END XNOR2x10_ASAP7_75t_SL

MACRO XNOR2x11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x11_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.292 0.504 4.048 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.476 0.252 3.816 0.324 ; 
        RECT 3.744 0.324 3.816 0.900 ; 
        RECT 0.828 0.900 3.816 0.972 ; 
    END 
  END Y
END XNOR2x11_ASAP7_75t_SL

MACRO XNOR2x12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x12_ASAP7_75t_SL 0 0 ; 
  SIZE 4.968 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 2.844 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 3.492 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 4.156 0.504 4.268 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.076 0.504 3.188 0.576 ; 
    END 
  END B
END XNOR2x12_ASAP7_75t_SL

MACRO XNOR2x14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x14_ASAP7_75t_SL 0 0 ; 
  SIZE 5.400 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 3.276 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 3.924 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 4.588 0.504 4.700 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.508 0.504 3.620 0.576 ; 
    END 
  END B
END XNOR2x14_ASAP7_75t_SL

MACRO XNOR2x16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x16_ASAP7_75t_SL 0 0 ; 
  SIZE 5.832 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 3.708 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 4.356 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 5.020 0.504 5.132 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.940 0.504 4.048 0.576 ; 
    END 
  END B
END XNOR2x16_ASAP7_75t_SL

MACRO XNOR2x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 1.892 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.324 1.548 0.396 ; 
        RECT 1.368 0.396 1.440 0.900 ; 
        RECT 0.828 0.900 1.548 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
END XNOR2x1_ASAP7_75t_SL

MACRO XNOR2x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 0.684 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 1.332 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.996 0.504 2.108 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END B
END XNOR2x2_ASAP7_75t_SL

MACRO XNOR2x4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x4_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 1.116 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 1.764 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.428 0.504 2.540 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.348 0.504 1.460 0.576 ; 
    END 
  END B
END XNOR2x4_ASAP7_75t_SL

MACRO XNOR2x5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x5_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.468 1.676 0.540 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XNOR2x5_ASAP7_75t_SL

MACRO XNOR2x7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x7_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.540 2.864 0.612 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.860 0.828 2.972 0.900 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
END XNOR2x7_ASAP7_75t_SL

MACRO XNOR2x9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x9_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.860 0.396 3.620 0.468 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.476 0.252 3.384 0.324 ; 
        RECT 3.312 0.324 3.384 0.900 ; 
        RECT 0.828 0.900 3.384 0.972 ; 
    END 
  END Y
END XNOR2x9_ASAP7_75t_SL

MACRO XOR2x10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x10_ASAP7_75t_SL 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 4.464 0.180 ; 
        RECT 4.392 0.180 4.464 0.900 ; 
        RECT 2.124 0.900 4.464 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x10_ASAP7_75t_SL

MACRO XOR2x11_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x11_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 4.048 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x11_ASAP7_75t_SL

MACRO XOR2x16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x16_ASAP7_75t_SL 0 0 ; 
  SIZE 5.832 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 5.760 0.180 ; 
        RECT 5.688 0.180 5.760 0.900 ; 
        RECT 2.124 0.900 5.760 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x16_ASAP7_75t_SL

MACRO XOR2x3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x3_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 2.324 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x3_ASAP7_75t_SL

MACRO XOR2x4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x4_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 3.168 0.180 ; 
        RECT 3.096 0.180 3.168 0.900 ; 
        RECT 2.124 0.900 3.168 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x4_ASAP7_75t_SL

MACRO XOR2x7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x7_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 3.188 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x7_ASAP7_75t_SL

MACRO XOR2x8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x8_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 4.032 0.180 ; 
        RECT 3.960 0.180 4.032 0.900 ; 
        RECT 2.124 0.900 4.032 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x8_ASAP7_75t_SL

MACRO XOR2x9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x9_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 3.620 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x9_ASAP7_75t_SL

MACRO INVx13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx13_ASAP7_75t_SL 0 0 ; 
  SIZE 3.240 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.168 0.180 ; 
        RECT 3.096 0.180 3.168 0.900 ; 
        RECT 0.396 0.900 3.168 0.972 ; 
    END 
  END Y
END INVx13_ASAP7_75t_SL

MACRO BUFx9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx9_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.980 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.980 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END A
END BUFx9_ASAP7_75t_SL

MACRO AND4x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND4x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
END AND4x1_ASAP7_75t_SL

MACRO OAI311xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI311xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B1
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C1
END OAI311xp33_ASAP7_75t_SL

MACRO OA222x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA222x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.288 0.396 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END A2
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B2
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END B1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END A1
END OA222x2_ASAP7_75t_SL

MACRO AND2x8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x8_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.872 0.180 ; 
        RECT 1.800 0.180 1.872 0.900 ; 
        RECT 0.396 0.900 1.872 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.496 2.304 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.444 2.088 0.636 ; 
    END 
  END A
END AND2x8_ASAP7_75t_SL

MACRO OA21x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21x2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.468 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A2
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B
END OA21x2_ASAP7_75t_SL

MACRO INVx15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx15_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.600 0.180 ; 
        RECT 3.528 0.180 3.600 0.900 ; 
        RECT 0.396 0.900 3.600 0.972 ; 
    END 
  END Y
END INVx15_ASAP7_75t_SL

MACRO AND2x10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x10_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.304 0.180 ; 
        RECT 2.232 0.180 2.304 0.900 ; 
        RECT 0.396 0.900 2.304 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.664 0.496 2.736 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.444 2.520 0.636 ; 
    END 
  END A
END AND2x10_ASAP7_75t_SL

MACRO AND2x16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x16_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 3.492 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 3.492 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.960 0.496 4.032 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.744 0.444 3.816 0.636 ; 
    END 
  END A
END AND2x16_ASAP7_75t_SL

MACRO BUFx13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx13_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 2.844 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 2.844 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.096 0.424 3.168 0.656 ; 
    END 
  END A
END BUFx13_ASAP7_75t_SL

MACRO DHLx8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx8_ASAP7_75t_SL 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.108 4.464 0.180 ; 
        RECT 4.392 0.180 4.464 0.900 ; 
        RECT 2.988 0.900 4.464 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx8_ASAP7_75t_SL

MACRO NAND5xp2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND5xp2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 1.116 0.972 ; 
    END 
  END Y
  PIN E
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END E
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
END NAND5xp2_ASAP7_75t_SL

MACRO AO333x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO333x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END C1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B3
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B1
  PIN C3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C3
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END C2
END AO333x1_ASAP7_75t_SL

MACRO OR2x16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x16_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.600 0.180 ; 
        RECT 3.528 0.180 3.600 0.900 ; 
        RECT 0.396 0.900 3.600 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.960 0.424 4.032 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.744 0.424 3.816 0.656 ; 
    END 
  END A
END OR2x16_ASAP7_75t_SL

MACRO OA22x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA22x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.288 0.396 0.360 0.756 ; 
        RECT 0.360 0.684 0.468 0.756 ; 
    END 
  END Y
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END B1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B2
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A2
END OA22x2_ASAP7_75t_SL

MACRO NAND4xp25_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp25_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.044 0.252 1.224 0.324 ; 
        RECT 1.152 0.324 1.224 0.900 ; 
        RECT 0.396 0.900 1.224 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END D
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C
END NAND4xp25_ASAP7_75t_SL

MACRO INVx4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx4_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.504 1.008 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.900 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 0.900 0.972 ; 
    END 
  END Y
END INVx4_ASAP7_75t_SL

MACRO DHLx4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx4_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.108 3.600 0.180 ; 
        RECT 3.528 0.180 3.600 0.900 ; 
        RECT 2.988 0.900 3.600 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx4_ASAP7_75t_SL

MACRO AND3x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B
END AND3x1_ASAP7_75t_SL

MACRO AND2x12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x12_ASAP7_75t_SL 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.736 0.180 ; 
        RECT 2.664 0.180 2.736 0.900 ; 
        RECT 0.396 0.900 2.736 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.096 0.496 3.168 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.880 0.444 2.952 0.636 ; 
    END 
  END A
END AND2x12_ASAP7_75t_SL

MACRO AO32x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO32x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.464 1.440 0.616 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.464 1.224 0.616 ; 
    END 
  END B1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.464 1.008 0.616 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.464 0.576 0.616 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.464 0.792 0.616 ; 
    END 
  END A2
END AO32x1_ASAP7_75t_SL

MACRO AO322x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO322x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.260 0.324 1.440 0.396 ; 
        RECT 1.368 0.396 1.440 0.684 ; 
        RECT 1.260 0.684 1.440 0.756 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END A2
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END B2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A3
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END B1
END AO322x2_ASAP7_75t_SL

MACRO INVx8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx8_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.504 1.656 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 1.764 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 1.764 0.972 ; 
    END 
  END Y
END INVx8_ASAP7_75t_SL

MACRO OAI332xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI332xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.692 0.252 2.088 0.324 ; 
        RECT 2.016 0.324 2.088 0.756 ; 
        RECT 0.828 0.756 2.088 0.828 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B3
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END C2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C1
END OAI332xp33_ASAP7_75t_SL

MACRO NOR2xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.252 0.792 0.324 ; 
        RECT 0.720 0.324 0.792 0.756 ; 
        RECT 0.612 0.756 0.792 0.828 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
END NOR2xp33_ASAP7_75t_SL

MACRO AO22x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO22x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A2
END AO22x1_ASAP7_75t_SL

MACRO DHLx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.324 0.252 0.756 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END CLK
END DHLx1_ASAP7_75t_SL

MACRO AND2x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.468 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A
END AND2x2_ASAP7_75t_SL

MACRO NAND3xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.080 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
END NAND3xp33_ASAP7_75t_SL

MACRO OR2x4_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x4_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.008 0.180 ; 
        RECT 0.936 0.180 1.008 0.900 ; 
        RECT 0.396 0.900 1.008 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A
END OR2x4_ASAP7_75t_SL

MACRO BUFx10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx10_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 2.196 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 2.196 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END A
END BUFx10_ASAP7_75t_SL

MACRO BUFx2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.080 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.288 0.396 0.360 0.972 ; 
        RECT 0.360 0.900 0.468 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A
END BUFx2_ASAP7_75t_SL

MACRO AOI321xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI321xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B2
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.828 0.108 1.656 0.180 ; 
        RECT 1.584 0.180 1.656 0.756 ; 
        RECT 1.260 0.756 1.656 0.828 ; 
    END 
  END Y
END AOI321xp33_ASAP7_75t_SL

MACRO AND5x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND5x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END D
  PIN E
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END E
END AND5x1_ASAP7_75t_SL

MACRO OAI222xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI222xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.692 0.252 2.088 0.324 ; 
        RECT 2.016 0.324 2.088 0.756 ; 
        RECT 0.612 0.756 2.088 0.828 ; 
    END 
  END Y
  PIN C2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C2
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END A2
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B1
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A1
END OAI222xp33_ASAP7_75t_SL

MACRO OR2x14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x14_ASAP7_75t_SL 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 3.168 0.180 ; 
        RECT 3.096 0.180 3.168 0.900 ; 
        RECT 0.396 0.900 3.168 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.528 0.424 3.600 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.424 3.384 0.656 ; 
    END 
  END A
END OR2x14_ASAP7_75t_SL

MACRO OR2x5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.116 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.116 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A
END OR2x5_ASAP7_75t_SL

MACRO OAI211xp5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI211xp5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.252 0.900 0.324 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END C
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
END OAI211xp5_ASAP7_75t_SL

MACRO AO21x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END B
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
END AO21x1_ASAP7_75t_SL

MACRO DFFLQNx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx1_ASAP7_75t_SL 0 0 ; 
  SIZE 4.320 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.484 0.360 0.596 ; 
    END 
  END CLK
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.484 1.224 0.596 ; 
    END 
  END D
  PIN QN
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.852 0.324 4.248 0.396 ; 
        RECT 4.176 0.396 4.248 0.684 ; 
        RECT 3.852 0.684 4.248 0.756 ; 
    END 
  END QN
END DFFLQNx1_ASAP7_75t_SL

MACRO NOR2x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 0.900 0.180 ; 
        RECT 0.504 0.180 0.576 0.684 ; 
        RECT 0.396 0.684 0.576 0.756 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END A
END NOR2x1_ASAP7_75t_SL

MACRO AND2x5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.116 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.116 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.496 1.656 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.444 1.440 0.636 ; 
    END 
  END A
END AND2x5_ASAP7_75t_SL

MACRO BUFx16_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx16_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 3.492 0.180 ; 
        RECT 0.288 0.180 0.360 0.972 ; 
        RECT 0.360 0.900 3.492 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.744 0.424 3.816 0.656 ; 
    END 
  END A
END BUFx16_ASAP7_75t_SL

MACRO INVx10_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx10_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 2.304 0.180 ; 
        RECT 2.232 0.180 2.304 0.900 ; 
        RECT 0.396 0.900 2.304 0.972 ; 
    END 
  END Y
END INVx10_ASAP7_75t_SL

MACRO OA331x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA331x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B2
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B3
  PIN C1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C1
END OA331x1_ASAP7_75t_SL

MACRO AO331x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO331x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A2
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A3
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A1
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B1
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END B2
  PIN B3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END B3
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END C
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.252 0.180 ; 
        RECT 0.072 0.180 0.144 0.756 ; 
        RECT 0.144 0.684 0.252 0.756 ; 
    END 
  END Y
END AO331x1_ASAP7_75t_SL

MACRO OR2x6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x6_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.440 0.180 ; 
        RECT 1.368 0.180 1.440 0.900 ; 
        RECT 0.396 0.900 1.440 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.424 1.656 0.656 ; 
    END 
  END A
END OR2x6_ASAP7_75t_SL

MACRO OAI221xp5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI221xp5_ASAP7_75t_SL 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.044 0.252 1.440 0.324 ; 
        RECT 1.368 0.324 1.440 0.900 ; 
        RECT 0.180 0.900 1.440 0.972 ; 
    END 
  END Y
  PIN B2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B2
  PIN B1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B1
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A1
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
END OAI221xp5_ASAP7_75t_SL

MACRO OA211x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA211x2_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.108 0.468 0.180 ; 
        RECT 0.288 0.180 0.360 0.756 ; 
        RECT 0.360 0.684 0.468 0.756 ; 
    END 
  END Y
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A2
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A1
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END C
END OA211x2_ASAP7_75t_SL

MACRO INVx7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx7_ASAP7_75t_SL 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.380 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.872 0.180 ; 
        RECT 1.800 0.180 1.872 0.900 ; 
        RECT 0.396 0.900 1.872 0.972 ; 
    END 
  END Y
END INVx7_ASAP7_75t_SL

MACRO AND2x15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x15_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 3.276 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 3.276 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.744 0.496 3.816 0.688 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.528 0.444 3.600 0.636 ; 
    END 
  END A
END AND2x15_ASAP7_75t_SL

MACRO DHLx7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx7_ASAP7_75t_SL 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.988 0.108 4.464 0.180 ; 
        RECT 4.392 0.180 4.464 0.900 ; 
        RECT 2.988 0.900 4.464 0.972 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END CLK
END DHLx7_ASAP7_75t_SL

MACRO AOI31xp33_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI31xp33_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.828 0.252 1.224 0.324 ; 
        RECT 1.152 0.324 1.224 0.756 ; 
        RECT 1.044 0.756 1.224 0.828 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END B
  PIN A1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END A1
  PIN A3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.424 0.360 0.656 ; 
    END 
  END A3
  PIN A2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2
END AOI31xp33_ASAP7_75t_SL

MACRO DLLx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.324 0.252 0.756 ; 
    END 
  END Q
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END CLK
END DLLx1_ASAP7_75t_SL

MACRO BUFx3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx3_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 0.684 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A
END BUFx3_ASAP7_75t_SL

MACRO BUFx7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx7_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.440 0.180 ; 
        RECT 1.368 0.180 1.440 0.900 ; 
        RECT 0.396 0.900 1.440 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.564 0.504 1.676 0.576 ; 
    END 
  END A
END BUFx7_ASAP7_75t_SL

MACRO OR2x7_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x7_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.548 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.548 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.800 0.424 1.872 0.656 ; 
    END 
  END A
END OR2x7_ASAP7_75t_SL

MACRO OR2x8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x8_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.396 0.108 1.872 0.180 ; 
        RECT 1.800 0.180 1.872 0.900 ; 
        RECT 0.396 0.900 1.872 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.016 0.424 2.088 0.656 ; 
    END 
  END A
END OR2x8_ASAP7_75t_SL

MACRO OR2x9_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x9_ASAP7_75t_SL 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.108 1.980 0.180 ; 
        RECT 0.072 0.180 0.144 0.972 ; 
        RECT 0.144 0.900 1.980 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.448 0.424 2.520 0.656 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 2.232 0.424 2.304 0.656 ; 
    END 
  END A
END OR2x9_ASAP7_75t_SL

MACRO OR3x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END A
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END C
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END B
END OR3x1_ASAP7_75t_SL

MACRO OR5x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR5x1_ASAP7_75t_SL 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.072 0.324 0.252 0.396 ; 
        RECT 0.072 0.396 0.144 0.972 ; 
        RECT 0.144 0.900 0.252 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.368 0.424 1.440 0.656 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END B
  PIN C
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.424 0.792 0.656 ; 
    END 
  END D
  PIN E
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END E
END OR5x1_ASAP7_75t_SL

MACRO SDFHx1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx1_ASAP7_75t_SL 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN SE
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.720 0.504 1.440 0.576 ; 
    END 
  END SE
  PIN D
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.484 0.360 0.596 ; 
    END 
  END D
  PIN CLK
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 3.312 0.484 3.384 0.596 ; 
    END 
  END CLK
  PIN SI
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.584 0.484 1.656 0.596 ; 
    END 
  END SI
  PIN QN
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 5.148 0.324 5.544 0.396 ; 
        RECT 5.472 0.396 5.544 0.684 ; 
        RECT 5.148 0.684 5.544 0.756 ; 
    END 
  END QN
END SDFHx1_ASAP7_75t_SL

MACRO XNOR2x13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x13_ASAP7_75t_SL 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.724 0.504 4.484 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.476 0.252 4.248 0.324 ; 
        RECT 4.176 0.324 4.248 0.900 ; 
        RECT 0.828 0.900 4.248 0.972 ; 
    END 
  END Y
END XNOR2x13_ASAP7_75t_SL

MACRO XNOR2x15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x15_ASAP7_75t_SL 0 0 ; 
  SIZE 5.184 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 4.156 0.504 4.916 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.476 0.252 4.680 0.324 ; 
        RECT 4.608 0.324 4.680 0.900 ; 
        RECT 0.828 0.900 4.680 0.972 ; 
    END 
  END Y
END XNOR2x15_ASAP7_75t_SL

MACRO XNOR2x3_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x3_ASAP7_75t_SL 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.564 0.504 2.324 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 1.476 0.252 2.088 0.324 ; 
        RECT 2.016 0.324 2.088 0.900 ; 
        RECT 0.828 0.900 2.088 0.972 ; 
    END 
  END Y
END XNOR2x3_ASAP7_75t_SL

MACRO XNOR2x6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x6_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 1.548 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 2.196 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.860 0.504 2.972 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.780 0.504 1.892 0.576 ; 
    END 
  END B
END XNOR2x6_ASAP7_75t_SL

MACRO XNOR2x8_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x8_ASAP7_75t_SL 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.180 0.108 1.980 0.180 ; 
        RECT 0.180 0.180 0.252 0.972 ; 
        RECT 0.252 0.900 2.628 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.292 0.504 3.404 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 2.212 0.504 2.324 0.576 ; 
    END 
  END B
END XNOR2x8_ASAP7_75t_SL

MACRO XOR2x12_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x12_ASAP7_75t_SL 0 0 ; 
  SIZE 4.968 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 4.896 0.180 ; 
        RECT 4.824 0.180 4.896 0.900 ; 
        RECT 2.124 0.900 4.896 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x12_ASAP7_75t_SL

MACRO XOR2x13_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x13_ASAP7_75t_SL 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 3.940 0.504 4.484 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x13_ASAP7_75t_SL

MACRO XOR2x14_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x14_ASAP7_75t_SL 0 0 ; 
  SIZE 5.400 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 5.328 0.180 ; 
        RECT 5.256 0.180 5.328 0.900 ; 
        RECT 2.124 0.900 5.328 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x14_ASAP7_75t_SL

MACRO XOR2x15_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x15_ASAP7_75t_SL 0 0 ; 
  SIZE 5.184 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 4.372 0.504 4.916 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x15_ASAP7_75t_SL

MACRO XOR2x1_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x1_ASAP7_75t_SL 0 0 ; 
  SIZE 2.160 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 1.892 0.576 ; 
    END 
  END A
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.828 0.108 1.548 0.180 ; 
        RECT 1.368 0.180 1.440 0.756 ; 
        RECT 1.440 0.684 1.548 0.756 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.288 0.324 0.792 0.396 ; 
        RECT 0.288 0.396 0.360 0.576 ; 
        RECT 0.720 0.396 0.792 0.576 ; 
    END 
  END B
END XOR2x1_ASAP7_75t_SL

MACRO XOR2x2_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x2_ASAP7_75t_SL 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.240 0.504 2.108 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.504 0.324 0.684 0.396 ; 
        RECT 0.504 0.396 0.576 0.972 ; 
        RECT 0.576 0.900 0.684 0.972 ; 
    END 
  END Y
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.268 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x2_ASAP7_75t_SL

MACRO XOR2x5_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x5_ASAP7_75t_SL 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 1.132 0.504 2.756 0.576 ; 
    END 
  END A
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.700 0.504 0.812 0.576 ; 
    END 
  END B
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal0 ;  
    END 
  END Y
END XOR2x5_ASAP7_75t_SL

MACRO XOR2x6_ASAP7_75t_SL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x6_ASAP7_75t_SL 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  PIN Y
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal1 ;  
        RECT 0.612 0.108 3.600 0.180 ; 
        RECT 3.528 0.180 3.600 0.900 ; 
        RECT 2.124 0.900 3.600 0.972 ; 
    END 
  END Y
  PIN B
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.484 0.504 0.596 0.576 ; 
    END 
  END B
  PIN A
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER metal2 ;  
        RECT 0.916 0.504 1.028 0.576 ; 
    END 
  END A
END XOR2x6_ASAP7_75t_SL

