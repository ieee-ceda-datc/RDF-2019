NangateOpenCellLibrary.mod.tech.lef