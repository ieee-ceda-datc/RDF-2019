VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS	2000 ;
END UNITS

MANUFACTURINGGRID	0.0025 ;

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  AREA 0.020000 ;
  WIDTH 0.065 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.072 ;
END VIA1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  AREA 0.020000 ;
  WIDTH 0.070 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.072 ;
END VIA2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  AREA 0.020000 ;
  WIDTH 0.070 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.072 ;
END VIA3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.072 ;
END VIA4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.072 ;
END VIA5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.072 ;
END VIA6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  AREA 0.020000 ;
  WIDTH 0.210 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal7

LAYER VIA7
  TYPE CUT ;
  SPACING 0.072 ;
END VIA7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.38 ;
  AREA 0.020000 ;
  WIDTH 0.210 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal8

LAYER VIA8
  TYPE CUT ;
  SPACING 0.072 ;
END VIA8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  AREA 0.020000 ;
  WIDTH 0.210 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal9

VIA VIA12 Default
  LAYER metal1 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA1 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal2 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12

VIA VIA23 Default
  LAYER metal2 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA2 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal3 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA23

VIA VIA34 Default
  LAYER metal3 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA3 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal4 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34

VIA VIA45 Default
  LAYER metal4 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA4 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal5 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA45

VIA VIA56 Default
  LAYER metal5 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA5 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal6 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA56

VIA VIA67 Default
  LAYER metal6 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA67

VIA VIA78 Default
  LAYER metal7 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal8 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA78

VIA VIA89 Default
  LAYER metal8 ;
	RECT -0.065000 -0.035000 0.065000 0.035000 ;
  LAYER VIA8 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal9 ;
	RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA89

END LIBRARY
