NangateOpenCellLibrary.mod.cell.lef