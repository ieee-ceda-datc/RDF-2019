NangateOpenCellLibrary.mod.lef